    Mac OS X            	   2   �      �                                      ATTR       �   �   "                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine E�a    I.    q/0081;00000000;; 