    Mac OS X            	   2   �      �                                      ATTR       �   �   "                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine Bf�c    d�    q/0081;00000000;; 