    Mac OS X            	   2   �      �                                      ATTR       �   �   "                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine �a    �>    q/0081;00000000;; 