LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY mux32to1 IS

    PORT (
        i_S : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
        i_D0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        i_D31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
        o_O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000");

END mux32to1;

ARCHITECTURE dataflow OF mux32to1 IS

BEGIN
    WITH i_S SELECT
        o_O <= i_D31 WHEN "11111",
        i_D30 WHEN "11110",
        i_D29 WHEN "11101",
        i_D28 WHEN "11100",
        i_D27 WHEN "11011",
        i_D26 WHEN "11010",
        i_D25 WHEN "11001",
        i_D24 WHEN "11000",
        i_D23 WHEN "10111",
        i_D22 WHEN "10110",
        i_D21 WHEN "10101",
        i_D20 WHEN "10100",
        i_D19 WHEN "10011",
        i_D18 WHEN "10010",
        i_D17 WHEN "10001",
        i_D16 WHEN "10000",
        i_D15 WHEN "01111",
        i_D14 WHEN "01110",
        i_D13 WHEN "01101",
        i_D12 WHEN "01100",
        i_D11 WHEN "01011",
        i_D10 WHEN "01010",
        i_D9 WHEN "01001",
        i_D8 WHEN "01000",
        i_D7 WHEN "00111",
        i_D6 WHEN "00110",
        i_D5 WHEN "00101",
        i_D4 WHEN "00100",
        i_D3 WHEN "00011",
        i_D2 WHEN "00010",
        i_D1 WHEN "00001",
        i_D0 WHEN "00000",
        "00000000000000000000000000000000" WHEN OTHERS;

END dataflow;